// Empty module for error testing
module empty_module(a, b, y);
  input logic a, b;
  output logic y;
endmodule
