// Assign statement test - OR
module assign_or(a, b, y);
  input logic a, b;
  output logic y;

  assign y = a | b;
endmodule
