// Assign statement test - AND
module assign_and(a, b, y);
  input logic a, b;
  output logic y;

  assign y = a & b;
endmodule
